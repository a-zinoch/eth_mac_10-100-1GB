`ifndef TIMESCALE
`define TIMESCALE

`timescale 1 ns / 100 ps

`endif //TIMESCALE