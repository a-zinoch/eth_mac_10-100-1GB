module CL_sync // syncronization Clocks by "Closed-loop"
	#(

	)(
		input clk_m
	, input clk_s
	,	input signal_i
	, input sig_ack_i


	);
endmodule
