module mem_contoller
	#(


	)(
			input 				reset_hard_i
		, input 				reset_i
		, input 				clk_i
		, input 				write_addr_cpu_tran
		, input 				write_addr_cpu_rec
		, input 				rec_OK
		, input [ 8:0 ]	





	)