`ifndef UNI_REG_PREDICTOR
`define UNI_REG_PREDICTOR

typedef uvm_reg_predictor#( sysbus_item ) uni_reg_predictor;

`endif //UNI_REG_PREDICTOR